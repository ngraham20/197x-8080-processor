----------------------------------------------------------
-- SEA_TOP
---------------------------------------------------------
library IEEE; 
use IEEE.STD_LOGIC_1164.all; 
use IEEE.STD_LOGIC_UNSIGNED.all;

entity sea_top is -- top-level design for testing
  port();
end;

---------------------------------------------------------
-- Architecture Definitions
---------------------------------------------------------

architecture sea_top of sea_top is

    end sea_top;
