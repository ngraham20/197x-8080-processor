----------------------------------------------------------
-- SEA_TOP
---------------------------------------------------------
library IEEE; 
use IEEE.STD_LOGIC_1164.all; 
use IEEE.STD_LOGIC_UNSIGNED.all;

entity sea_top is -- top-level design for testing
  port();
end;

---------------------------------------------------------
-- Architecture Definitions
---------------------------------------------------------

architecture sea_top of sea_top is

    end sea_top;
    
    
-- TODO finish the top
-- TODO finish the CU
-- TODO fix the srr and srl errors in the alu
-- TODO bit stuff
-- TODO bug fixes
-- TODO create test sea program
